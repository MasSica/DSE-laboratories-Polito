LIBRARY ieee;USE ieee.std_logic_1164.all; USE ieee.numeric_std.all;entity stage_one is PORT (add,badd : in std_logic_vector(3 downto 0);cin: in std_logic;sum: out std_logic_vector(3 downto 0);cout: out std_logic);end stage_one;architecture behavior of stage_one is signal carry: std_logic_vector(2 downto 0);component full_add is PORT (a,b: in std_logic;      c_in: in std_logic;      c_out,s: out std_logic);end component;begin fa1:full_add PORT MAP(add(0),badd(0),'0',carry(0),sum(0));fa2:full_add PORT MAP(add(1),badd(1),carry(0),carry(1),sum(1));fa3:full_add PORT MAP(add(2),badd(2),carry(1),carry(2),sum(2));fa4:full_add PORT MAP(add(3),badd(3),carry(2),cout,sum(3));end behavior;
LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.numeric_std.all;ENTITY reaction_tb ISEND reaction_tb;ARCHITECTURE arch of reaction_tb issignal sw_tb: unsigned(7 downto 0);	signal clock_tb: std_logic;signal KEY0_tb,KEY3_tb: std_logic;signal LEDR0_tb: std_logic;signal HEX3_tb,HEX2_tb,HEX1_tb,HEX0_tb:std_logic_vector(0 to 6);component reaction isport( SW: in unsigned (7 downto 0);clock_50: in std_logic;KEY0,KEY3:in std_logic;LEDR0: out std_logic;HEX3,HEX2,HEX1,HEX0:out std_logic_vector(0 to 6));end component;BEGINuut: reaction PORT MAP(sw_tb,clock_tb,KEY0_tb,KEY3_tb,LEDR0_tb,HEX3_tb,HEX2_tb,HEX1_tb,HEX0_tb);processbeginsw_tb <= "00000010";KEY0_tb<='1';wait for 25 ns;KEY0_tb<='0';wait for 1500 ns;KEY3_tb<='1';wait for 25 ns;KEY3_tb<='0';wait for 500 ns;KEY0_tb<='1';wait for 25 ns;KEY0_tb<='0';wait for 2000 ns;KEY3_tb<='1';wait for 25 ns;KEY3_tb<='0';wait;end process;PROCESS(clock_tb) BEGINif clock_tb='U' then	clock_tb<='0' after 10 ns;else	clock_tb<= not clock_tb after 10 ns;end if;end process;END arch;